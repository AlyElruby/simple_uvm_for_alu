package alu_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "alu_transaction.svh"
    `include "alu_sequencer.svh"
    `include "alu_scoreboard.svh"
    `include "alu_driver.svh"
    `include "alu_monitor.svh"
    `include "alu_agent.svh"
    `include "alu_env.svh"
    `include "alu_test.svh"
endpackage